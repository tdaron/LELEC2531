module modulo();
endmodule;
